module moduleName (
    input wire, 
    output wire
);
    
endmodule